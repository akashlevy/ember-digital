
//^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^
// GF(5)
//^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^

function automatic [9:0] fn_bch_dec_gf5;
input[30:0] d;

reg [9:0] p;
begin

p[0] = d[0]^ d[1]^ d[3]^ d[5]^ d[7]^ d[8]^ d[9]^ d[10]^ d[13]^ d[16]^ d[18]^ d[21];
p[1] = d[1]^ d[2]^ d[4]^ d[6]^ d[8]^ d[9]^ d[10]^ d[11]^ d[14]^ d[17]^ d[19]^ d[22];
p[2] = d[2]^ d[3]^ d[5]^ d[7]^ d[9]^ d[10]^ d[11]^ d[12]^ d[15]^ d[18]^ d[20]^ d[23];
p[3] = d[0]^ d[1]^ d[4]^ d[5]^ d[6]^ d[7]^ d[9]^ d[11]^ d[12]^ d[18]^ d[19]^ d[24];
p[4] = d[1]^ d[2]^ d[5]^ d[6]^ d[7]^ d[8]^ d[10]^ d[12]^ d[13]^ d[19]^ d[20]^ d[25];
p[5] = d[0]^ d[1]^ d[2]^ d[5]^ d[6]^ d[10]^ d[11]^ d[14]^	d[16]^ d[18]^ d[20]^ d[26];
p[6] = d[0]^ d[2]^ d[5]^ d[6]^ d[8]^ d[9]^ d[10]^ d[11]^ d[12]^ d[13]^ d[15]^ d[16]^ d[17]^ d[18]^ d[19]^ d[27];
p[7] = d[1]^ d[3]^ d[6]^ d[7]^ d[9]^ d[10]^ d[11]^ d[12]^ d[13]^ d[14]^ d[16]^ d[17]^ d[18]^ d[19]^ d[20]^ d[28];
p[8] = d[0]^ d[1]^ d[2]^ d[3]^ d[4]^ d[5]^ d[9]^ d[11]^ d[12]^ d[14]^ d[15]^	d[16]^ d[17]^ d[19]^ d[20]^ d[29];
p[9] = d[0]^ d[2]^ d[4]^ d[6]^ d[7]^ d[8]^ d[9]^ d[12]^ d[15]^	d[17]^ d[20]^ d[30];

fn_bch_dec_gf5 = p;
end	

endfunction // fn_bch_dec_gf5

